module top_module (
  output out
);
  assign out = 1'b0; // 输出固定为0的信号
endmodule
