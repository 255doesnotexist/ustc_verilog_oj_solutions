module top_module (
  output out
);
  assign out = 1'b1; // 输出固定为1的信号
endmodule
