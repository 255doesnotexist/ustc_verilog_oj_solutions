module top_module( input in, output out );
// 请用户在下方编辑代码
  assign out = !in;
//用户编辑到此为止
endmodule