module top_module( 
    input a,b,c,
    output w,x,y,z );
// 请用户在下方编辑代码
    assign a_wire = a;
    assign b_wire = b;
    assign c_wire = c;

    assign w = a_wire;
    assign x = b_wire;
    assign y = b_wire;
    assign z = c_wire;
//用户编辑到此为止
endmodule
